`include "spi_master_slave_rtl.v"
`include "top.v"
`include "transac.sv"
`include "intf.sv"
`include "gen.sv"
`include "drv.sv"
`include "mon.sv"
`include "scb.sv"
`include "tb.sv"
